// Verilog netlist created by Tang Dynasty v5.9.122301
// Sun Dec  1 11:04:47 2024

`timescale 1ns / 1ps
module top_CIC_0
  (
  clk,
  din,
  din_en,
  rst,
  dout,
  dout_en
  );

  input clk;
  input [15:0] din;
  input din_en;
  input rst;
  output [28:0] dout;
  output dout_en;

  wire [2:0] al_1deac949;
  wire [3:0] al_54f1bd90;
  wire [28:0] al_eb2ab31;
  wire [28:0] al_480f15b7;
  wire [28:0] al_8f688f54;
  wire [28:0] al_e9628d6d;
  wire [28:0] al_4fe8581e;
  wire [28:0] al_6d487ee0;
  wire [28:0] al_7d3eb7bc;
  wire [28:0] al_feb3b069;
  wire [28:0] al_2c916a43;
  wire [28:0] al_be8c6636;
  wire [28:0] al_62f4aab;
  wire [28:0] al_5414e669;
  wire [28:0] al_4e1fa175;
  wire [28:0] al_cd893e44;
  wire [28:0] al_b27b90b2;
  wire [28:0] al_4873fb93;
  wire [28:0] al_9955f70;
  wire [28:0] al_14ec71c5;
  wire [28:0] al_d9b93292;
  wire [28:0] al_afdc4416;
  wire [28:0] al_5e11d7be;
  wire [28:0] al_1d216208;
  wire [28:0] al_6d689829;
  wire [28:0] al_1358e4cb;
  wire [28:0] al_ac1e65eb;
  wire al_5fed0cdc;
  wire al_2eeaca0f;
  wire al_711addca;
  wire al_317aa4ea;
  wire al_58f3b920;
  wire al_d6bc4586;
  wire al_3ce59305;
  wire al_700a31d9;
  wire al_53dc503e;
  wire al_277f2230;
  wire al_e4916434;
  wire al_3c6b44d0;
  wire al_210843f4;
  wire al_f6f3ead6;
  wire al_6ce64f20;
  wire al_25624ff1;
  wire al_27e555a3;
  wire al_7a35791a;
  wire al_994b351d;
  wire al_5f5bdd6f;
  wire al_423e8511;
  wire al_5dd3996b;
  wire al_1d1e96a3;
  wire al_93780002;
  wire al_3230880;
  wire al_881729c4;
  wire al_761c35be;
  wire al_7d4513e7;
  wire al_7b7f1ce4;
  wire al_e3df519b;
  wire al_44f5ebdc;
  wire al_a05a0af7;
  wire al_87331174;
  wire al_e6ce6c9f;
  wire al_4d39c51c;
  wire al_77098fec;
  wire al_f7b6239e;
  wire al_4100520;
  wire al_9980245b;
  wire al_2a38127a;
  wire al_32930761;
  wire al_335dce21;
  wire al_3e9c55c9;
  wire al_b1b1fd25;
  wire al_c0541eeb;
  wire al_8fa663c7;
  wire al_aea9f159;
  wire al_b5999e8a;
  wire al_4e02a214;
  wire al_e4bb6517;
  wire al_c7d5f7d9;
  wire al_aa0a4406;
  wire al_2936d63e;
  wire al_c33532a1;
  wire al_a1d7e557;
  wire al_535bcb2a;
  wire al_8e96be84;
  wire al_7f24ef3b;
  wire al_ea32c6e1;
  wire al_2ac97405;
  wire al_a0ebd25;
  wire al_f77a35ee;
  wire al_2902a00c;
  wire al_94925fa9;
  wire al_51a70210;
  wire al_fbeca432;
  wire al_ca5b12bc;
  wire al_b49c276a;
  wire al_a23af5a4;
  wire al_fe2986b6;
  wire al_875c79d9;
  wire al_d21ff3d4;
  wire al_20da7cd1;
  wire al_4b6c2990;
  wire al_2a9315a6;
  wire al_b9c5d958;
  wire al_56630a35;
  wire al_a1b0b17a;
  wire al_7b07bb65;
  wire al_9df2af8f;
  wire al_df20ca5b;
  wire al_ab6a0e7;
  wire al_3f047599;
  wire al_b4d1b2a2;
  wire al_469cb985;
  wire al_ffb568cb;
  wire al_8f0bd67f;
  wire al_b0d09b8;
  wire al_94c23594;
  wire al_d203b819;
  wire al_c5f97e65;
  wire al_5aa7ca6a;
  wire al_c709f85a;
  wire al_26a0aae;
  wire al_94b1300d;
  wire al_1e9cae1d;
  wire al_13006735;
  wire al_bbd9355;
  wire al_8f481ef9;
  wire al_9ab66270;
  wire al_4dcb26fa;
  wire al_d0181d13;
  wire al_b08aad73;
  wire al_c1c08587;
  wire al_689cec14;
  wire al_9ddddc8e;
  wire al_41a92fc7;
  wire al_d4d70e4b;
  wire al_e800c9ef;
  wire al_5cf39772;
  wire al_339b3bc;
  wire al_c6da537;
  wire al_35361f12;
  wire al_c6028b1e;
  wire al_87b345e3;
  wire al_29505f4f;
  wire al_aa8f2cd8;
  wire al_685d248f;
  wire al_cfde68ec;
  wire al_5c1d9288;
  wire al_1f7974b0;
  wire al_c964d6b6;
  wire al_d5344387;
  wire al_944a7435;
  wire al_16b99b31;
  wire al_5c3c8bc3;
  wire al_83d3841d;
  wire al_21712447;
  wire al_e26baa7c;
  wire al_bd632267;
  wire al_7b0a2fb3;
  wire al_b8ace6d9;
  wire al_18580a3b;
  wire al_830367be;
  wire al_92e30c9d;
  wire al_6566c57e;
  wire al_29ad0e3a;
  wire al_51513f80;
  wire al_1cd5a819;
  wire al_11e537d;
  wire al_5d5b70cd;
  wire al_397e2eb4;
  wire al_60062243;
  wire al_14a9163b;
  wire al_ca0bd035;
  wire al_10ad2d4;
  wire al_4b7e6f4c;
  wire al_dc48d934;
  wire al_65f78d31;
  wire al_9f58115d;
  wire al_6678a2d9;
  wire al_d662cc5f;
  wire al_121b0ac0;
  wire al_74c02a6e;
  wire al_2c19a30d;
  wire al_30e98b36;
  wire al_dff2b81e;
  wire al_7e683184;
  wire al_b5ad59ae;
  wire al_fdc784df;
  wire al_8625eee6;
  wire al_b46339ca;
  wire al_47553d9c;
  wire al_e55eeb92;
  wire al_2bd76071;
  wire al_f5c68653;
  wire al_7b6818a7;
  wire al_ce1229f8;
  wire al_77221701;
  wire al_c6a9c727;
  wire al_e5f7a519;
  wire al_c65e25f4;
  wire al_a839234c;
  wire al_e0116105;
  wire al_b7706566;
  wire al_32713696;
  wire al_58c1d211;
  wire al_f6e6833c;
  wire al_d6b08360;
  wire al_ab39c04d;
  wire al_a1a76be0;
  wire al_80b80f4;
  wire al_a8099213;
  wire al_89797e8b;
  wire al_d4fb750d;
  wire al_c0a4beaf;
  wire al_f1885c7b;
  wire al_406fb43d;
  wire al_2ae006a6;
  wire al_25a1ab81;
  wire al_7bc6bbc7;
  wire al_5d510d59;
  wire al_d82381d;
  wire al_9f37eb9f;
  wire al_3fca7;
  wire al_22c2b9e6;
  wire al_72694321;
  wire al_5e0efc9d;
  wire al_4218870a;
  wire al_debafe7e;
  wire al_fd1c7e35;
  wire al_f4a4c863;
  wire al_47aec73d;
  wire al_da97260d;
  wire al_54f6d4d2;
  wire al_ca0ec285;
  wire al_8a5edc6c;
  wire al_82b795a6;
  wire al_cb347ae8;
  wire al_fbe9b8eb;
  wire al_855a8144;
  wire al_50dcf253;
  wire al_5a7c92db;
  wire al_12f77c35;
  wire al_c2eaa9c5;
  wire al_7c0b757b;
  wire al_3ec6aa29;
  wire al_3048204c;
  wire al_105495bd;
  wire al_3b6a1fd8;
  wire al_7025ee8e;
  wire al_d397fa50;
  wire al_e1210075;
  wire al_6fdacc18;
  wire al_9dd79649;
  wire al_9e87a365;
  wire al_ff6a88f6;
  wire al_404f5287;
  wire al_5d53cef6;
  wire al_4ed44021;
  wire al_f392c8e6;
  wire al_cc8f42a5;
  wire al_3c97da5f;
  wire al_3bce7a34;
  wire al_418f7602;
  wire al_dd04a5ca;
  wire al_461ca1b0;
  wire al_dec8e5a2;
  wire al_66eadc2c;
  wire al_60c7c36e;
  wire al_8f3aa2df;
  wire al_fb131175;
  wire al_90fed4e7;
  wire al_10238dc7;
  wire al_8b4171c8;
  wire al_2c346a44;
  wire al_36624d30;
  wire al_438b278b;
  wire al_de0bda5;
  wire al_89db50f8;
  wire al_d2835c11;
  wire al_e0e4e676;
  wire al_685ac330;
  wire al_bc1a95db;
  wire al_c7938c90;
  wire al_3b1bd3d;
  wire al_1c7d78dc;
  wire al_c4c4b744;
  wire al_82fc816d;
  wire al_85782b8c;
  wire al_52d5f2ec;
  wire al_ce46c960;
  wire al_8d67c17b;
  wire al_6b121a3b;
  wire al_2867582b;
  wire al_62124ca0;
  wire al_2e19f2fe;
  wire al_a1734311;
  wire al_9b8ea422;
  wire al_d548edf7;
  wire al_6bb3744a;
  wire al_70d5777e;
  wire al_31957fb7;
  wire al_40f92736;
  wire al_bc0758d;
  wire al_98711f8a;
  wire al_62e158f1;
  wire al_bd8fc407;
  wire al_b1815462;
  wire al_e23d25b3;
  wire al_62be7f6f;
  wire al_58af7ea5;
  wire al_6b633f05;
  wire al_fcebab7e;
  wire al_53c60bff;
  wire al_1b2cf291;
  wire al_e060e572;
  wire al_d57ca002;
  wire al_9f2e787e;
  wire al_560a769;
  wire al_f76ae046;
  wire al_1b884b48;
  wire al_45855c0b;
  wire al_3a284b58;
  wire al_8b833a2e;
  wire al_65b98507;
  wire al_3fe5f260;
  wire al_81c141dd;
  wire al_fd840f8c;
  wire al_4705248d;
  wire al_229e7e2c;

  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_2d21f01f (
    .a(1'b0),
    .o({al_5fed0cdc,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8fdb2b60 (
    .a(al_eb2ab31[0]),
    .b(din[0]),
    .c(al_5fed0cdc),
    .o({al_2eeaca0f,al_480f15b7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_24d032cc (
    .a(al_eb2ab31[1]),
    .b(din[1]),
    .c(al_2eeaca0f),
    .o({al_711addca,al_480f15b7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_19519ce (
    .a(al_eb2ab31[2]),
    .b(din[2]),
    .c(al_711addca),
    .o({al_317aa4ea,al_480f15b7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_df4222bb (
    .a(al_eb2ab31[3]),
    .b(din[3]),
    .c(al_317aa4ea),
    .o({al_58f3b920,al_480f15b7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a2e63e7a (
    .a(al_eb2ab31[4]),
    .b(din[4]),
    .c(al_58f3b920),
    .o({al_d6bc4586,al_480f15b7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a546e215 (
    .a(al_eb2ab31[5]),
    .b(din[5]),
    .c(al_d6bc4586),
    .o({al_3ce59305,al_480f15b7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e4833917 (
    .a(al_eb2ab31[6]),
    .b(din[6]),
    .c(al_3ce59305),
    .o({al_700a31d9,al_480f15b7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_204285ef (
    .a(al_eb2ab31[7]),
    .b(din[7]),
    .c(al_700a31d9),
    .o({al_53dc503e,al_480f15b7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7ea63a6f (
    .a(al_eb2ab31[8]),
    .b(din[8]),
    .c(al_53dc503e),
    .o({al_277f2230,al_480f15b7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_77257231 (
    .a(al_eb2ab31[9]),
    .b(din[9]),
    .c(al_277f2230),
    .o({al_e4916434,al_480f15b7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bc5eb54d (
    .a(al_eb2ab31[10]),
    .b(din[10]),
    .c(al_e4916434),
    .o({al_3c6b44d0,al_480f15b7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2d23a90d (
    .a(al_eb2ab31[11]),
    .b(din[11]),
    .c(al_3c6b44d0),
    .o({al_210843f4,al_480f15b7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_de47ac8e (
    .a(al_eb2ab31[12]),
    .b(din[12]),
    .c(al_210843f4),
    .o({al_f6f3ead6,al_480f15b7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c889a44a (
    .a(al_eb2ab31[13]),
    .b(din[13]),
    .c(al_f6f3ead6),
    .o({al_6ce64f20,al_480f15b7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_77d22e77 (
    .a(al_eb2ab31[14]),
    .b(din[14]),
    .c(al_6ce64f20),
    .o({al_25624ff1,al_480f15b7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f506b27d (
    .a(al_eb2ab31[15]),
    .b(din[15]),
    .c(al_25624ff1),
    .o({al_27e555a3,al_480f15b7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_30a8497b (
    .a(al_eb2ab31[16]),
    .b(din[15]),
    .c(al_27e555a3),
    .o({al_7a35791a,al_480f15b7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_32d88032 (
    .a(al_eb2ab31[17]),
    .b(din[15]),
    .c(al_7a35791a),
    .o({al_994b351d,al_480f15b7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6862943f (
    .a(al_eb2ab31[18]),
    .b(din[15]),
    .c(al_994b351d),
    .o({al_5f5bdd6f,al_480f15b7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_31eb4985 (
    .a(al_eb2ab31[19]),
    .b(din[15]),
    .c(al_5f5bdd6f),
    .o({al_423e8511,al_480f15b7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cd217c4a (
    .a(al_eb2ab31[20]),
    .b(din[15]),
    .c(al_423e8511),
    .o({al_5dd3996b,al_480f15b7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a707256f (
    .a(al_eb2ab31[21]),
    .b(din[15]),
    .c(al_5dd3996b),
    .o({al_1d1e96a3,al_480f15b7[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_92580e69 (
    .a(al_eb2ab31[22]),
    .b(din[15]),
    .c(al_1d1e96a3),
    .o({al_93780002,al_480f15b7[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ee343458 (
    .a(al_eb2ab31[23]),
    .b(din[15]),
    .c(al_93780002),
    .o({al_3230880,al_480f15b7[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_556ce633 (
    .a(al_eb2ab31[24]),
    .b(din[15]),
    .c(al_3230880),
    .o({al_881729c4,al_480f15b7[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_aefd8b68 (
    .a(al_eb2ab31[25]),
    .b(din[15]),
    .c(al_881729c4),
    .o({al_761c35be,al_480f15b7[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_32ed25d3 (
    .a(al_eb2ab31[26]),
    .b(din[15]),
    .c(al_761c35be),
    .o({al_7d4513e7,al_480f15b7[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2fcc6939 (
    .a(al_eb2ab31[27]),
    .b(din[15]),
    .c(al_7d4513e7),
    .o({al_7b7f1ce4,al_480f15b7[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d39fb125 (
    .a(al_eb2ab31[28]),
    .b(din[15]),
    .c(al_7b7f1ce4),
    .o({open_n3,al_480f15b7[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_6c65e6ec (
    .a(1'b0),
    .o({al_e3df519b,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7a814cc1 (
    .a(al_2c916a43[8]),
    .b(al_7d3eb7bc[8]),
    .c(al_4100520),
    .o({al_9980245b,al_be8c6636[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f0f1414 (
    .a(al_2c916a43[9]),
    .b(al_7d3eb7bc[9]),
    .c(al_9980245b),
    .o({al_2a38127a,al_be8c6636[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bd625e74 (
    .a(al_2c916a43[10]),
    .b(al_7d3eb7bc[10]),
    .c(al_2a38127a),
    .o({al_32930761,al_be8c6636[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f66cc420 (
    .a(al_2c916a43[11]),
    .b(al_7d3eb7bc[11]),
    .c(al_32930761),
    .o({al_335dce21,al_be8c6636[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_be113f82 (
    .a(al_2c916a43[12]),
    .b(al_7d3eb7bc[12]),
    .c(al_335dce21),
    .o({al_3e9c55c9,al_be8c6636[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_197ca113 (
    .a(al_2c916a43[13]),
    .b(al_7d3eb7bc[13]),
    .c(al_3e9c55c9),
    .o({al_b1b1fd25,al_be8c6636[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_16c07b12 (
    .a(al_2c916a43[14]),
    .b(al_7d3eb7bc[14]),
    .c(al_b1b1fd25),
    .o({al_c0541eeb,al_be8c6636[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e77d29a3 (
    .a(al_2c916a43[15]),
    .b(al_7d3eb7bc[15]),
    .c(al_c0541eeb),
    .o({al_8fa663c7,al_be8c6636[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a710bda1 (
    .a(al_2c916a43[16]),
    .b(al_7d3eb7bc[16]),
    .c(al_8fa663c7),
    .o({al_aea9f159,al_be8c6636[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_21783b3a (
    .a(al_2c916a43[17]),
    .b(al_7d3eb7bc[17]),
    .c(al_aea9f159),
    .o({al_b5999e8a,al_be8c6636[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c2cd2d4e (
    .a(al_2c916a43[0]),
    .b(al_7d3eb7bc[0]),
    .c(al_e3df519b),
    .o({al_44f5ebdc,al_be8c6636[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7bffdcb2 (
    .a(al_2c916a43[18]),
    .b(al_7d3eb7bc[18]),
    .c(al_b5999e8a),
    .o({al_4e02a214,al_be8c6636[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_11f7f27b (
    .a(al_2c916a43[19]),
    .b(al_7d3eb7bc[19]),
    .c(al_4e02a214),
    .o({al_e4bb6517,al_be8c6636[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_791e3201 (
    .a(al_2c916a43[20]),
    .b(al_7d3eb7bc[20]),
    .c(al_e4bb6517),
    .o({al_c7d5f7d9,al_be8c6636[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c98cb61e (
    .a(al_2c916a43[21]),
    .b(al_7d3eb7bc[21]),
    .c(al_c7d5f7d9),
    .o({al_aa0a4406,al_be8c6636[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e40ddbb4 (
    .a(al_2c916a43[22]),
    .b(al_7d3eb7bc[22]),
    .c(al_aa0a4406),
    .o({al_2936d63e,al_be8c6636[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a6dbf441 (
    .a(al_2c916a43[23]),
    .b(al_7d3eb7bc[23]),
    .c(al_2936d63e),
    .o({al_c33532a1,al_be8c6636[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2fa277d8 (
    .a(al_2c916a43[24]),
    .b(al_7d3eb7bc[24]),
    .c(al_c33532a1),
    .o({al_a1d7e557,al_be8c6636[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5b9299c0 (
    .a(al_2c916a43[25]),
    .b(al_7d3eb7bc[25]),
    .c(al_a1d7e557),
    .o({al_535bcb2a,al_be8c6636[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6a0b44d (
    .a(al_2c916a43[26]),
    .b(al_7d3eb7bc[26]),
    .c(al_535bcb2a),
    .o({al_8e96be84,al_be8c6636[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6a1f217 (
    .a(al_2c916a43[27]),
    .b(al_7d3eb7bc[27]),
    .c(al_8e96be84),
    .o({al_7f24ef3b,al_be8c6636[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_39375266 (
    .a(al_2c916a43[1]),
    .b(al_7d3eb7bc[1]),
    .c(al_44f5ebdc),
    .o({al_a05a0af7,al_be8c6636[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_57fd69b4 (
    .a(al_2c916a43[28]),
    .b(al_7d3eb7bc[28]),
    .c(al_7f24ef3b),
    .o({open_n7,al_be8c6636[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1be482f2 (
    .a(al_2c916a43[2]),
    .b(al_7d3eb7bc[2]),
    .c(al_a05a0af7),
    .o({al_87331174,al_be8c6636[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_63d33a4b (
    .a(al_2c916a43[3]),
    .b(al_7d3eb7bc[3]),
    .c(al_87331174),
    .o({al_e6ce6c9f,al_be8c6636[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c797f8a4 (
    .a(al_2c916a43[4]),
    .b(al_7d3eb7bc[4]),
    .c(al_e6ce6c9f),
    .o({al_4d39c51c,al_be8c6636[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7f656e5 (
    .a(al_2c916a43[5]),
    .b(al_7d3eb7bc[5]),
    .c(al_4d39c51c),
    .o({al_77098fec,al_be8c6636[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b11b3677 (
    .a(al_2c916a43[6]),
    .b(al_7d3eb7bc[6]),
    .c(al_77098fec),
    .o({al_f7b6239e,al_be8c6636[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f1a11535 (
    .a(al_2c916a43[7]),
    .b(al_7d3eb7bc[7]),
    .c(al_f7b6239e),
    .o({al_4100520,al_be8c6636[7]}));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_d0c3c85e (
    .a(al_1deac949[0]),
    .o(al_da97260d));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+~(A)*B*C)"),
    .INIT(8'h46))
    al_90fbe134 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .c(al_1deac949[2]),
    .o(al_54f1bd90[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+~(A)*~(B)*C+~(A)*B*C)"),
    .INIT(8'h58))
    al_68639997 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .c(al_1deac949[2]),
    .o(al_54f1bd90[2]));
  AL_DFF_X al_eb711602 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_da97260d),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_X al_8e369bed (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_54f1bd90[1]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_X al_ace4f707 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_54f1bd90[2]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_X al_a83b24f5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_229e7e2c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout_en));
  AL_DFF_X al_5791a65c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[0]));
  AL_DFF_X al_8efda135 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[9]));
  AL_DFF_X al_61567a29 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[10]));
  AL_DFF_X al_ca0d43a5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[11]));
  AL_DFF_X al_b736491a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[12]));
  AL_DFF_X al_c86a1a3b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[13]));
  AL_DFF_X al_7dc951b7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[14]));
  AL_DFF_X al_391c3fe4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[15]));
  AL_DFF_X al_3c09d507 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[16]));
  AL_DFF_X al_a9cf0690 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[17]));
  AL_DFF_X al_85625e02 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[18]));
  AL_DFF_X al_eab0872a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[1]));
  AL_DFF_X al_cb822b6f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[19]));
  AL_DFF_X al_98310e40 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[20]));
  AL_DFF_X al_57ac6c81 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[21]));
  AL_DFF_X al_49a1b852 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[22]));
  AL_DFF_X al_b5bb55fc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[23]));
  AL_DFF_X al_295aa775 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[24]));
  AL_DFF_X al_b79d4840 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[25]));
  AL_DFF_X al_7fe3aaf6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[26]));
  AL_DFF_X al_284e7e34 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[27]));
  AL_DFF_X al_bebccd1b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[28]));
  AL_DFF_X al_b70fcc76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[2]));
  AL_DFF_X al_75019a17 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[3]));
  AL_DFF_X al_798d38ff (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[4]));
  AL_DFF_X al_22266b1a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[5]));
  AL_DFF_X al_c7ee36c5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[6]));
  AL_DFF_X al_c4eed9ba (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[7]));
  AL_DFF_X al_5f3179e4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1358e4cb[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(dout[8]));
  AL_DFF_X al_de6e4cf3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(din_en),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_54f6d4d2));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fce83d32 (
    .a(al_eb2ab31[7]),
    .b(al_8f688f54[7]),
    .c(al_5a7c92db),
    .o({al_12f77c35,al_e9628d6d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dd2124b4 (
    .a(al_eb2ab31[8]),
    .b(al_8f688f54[8]),
    .c(al_12f77c35),
    .o({al_c2eaa9c5,al_e9628d6d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec563035 (
    .a(al_eb2ab31[9]),
    .b(al_8f688f54[9]),
    .c(al_c2eaa9c5),
    .o({al_7c0b757b,al_e9628d6d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f4d2e6b5 (
    .a(al_eb2ab31[10]),
    .b(al_8f688f54[10]),
    .c(al_7c0b757b),
    .o({al_3ec6aa29,al_e9628d6d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b48d723f (
    .a(al_eb2ab31[11]),
    .b(al_8f688f54[11]),
    .c(al_3ec6aa29),
    .o({al_3048204c,al_e9628d6d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bcb6bfa3 (
    .a(al_eb2ab31[12]),
    .b(al_8f688f54[12]),
    .c(al_3048204c),
    .o({al_105495bd,al_e9628d6d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f73d1c0c (
    .a(al_eb2ab31[13]),
    .b(al_8f688f54[13]),
    .c(al_105495bd),
    .o({al_3b6a1fd8,al_e9628d6d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c670403a (
    .a(al_eb2ab31[14]),
    .b(al_8f688f54[14]),
    .c(al_3b6a1fd8),
    .o({al_7025ee8e,al_e9628d6d[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_be53845b (
    .a(al_eb2ab31[15]),
    .b(al_8f688f54[15]),
    .c(al_7025ee8e),
    .o({al_d397fa50,al_e9628d6d[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_586da07d (
    .a(al_eb2ab31[16]),
    .b(al_8f688f54[16]),
    .c(al_d397fa50),
    .o({al_e1210075,al_e9628d6d[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_28d1cd6 (
    .a(1'b0),
    .o({al_ca0ec285,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f74e7eb (
    .a(al_eb2ab31[17]),
    .b(al_8f688f54[17]),
    .c(al_e1210075),
    .o({al_6fdacc18,al_e9628d6d[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f544a4d7 (
    .a(al_eb2ab31[18]),
    .b(al_8f688f54[18]),
    .c(al_6fdacc18),
    .o({al_9dd79649,al_e9628d6d[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_39814d66 (
    .a(al_eb2ab31[19]),
    .b(al_8f688f54[19]),
    .c(al_9dd79649),
    .o({al_9e87a365,al_e9628d6d[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_acc18a81 (
    .a(al_eb2ab31[20]),
    .b(al_8f688f54[20]),
    .c(al_9e87a365),
    .o({al_ff6a88f6,al_e9628d6d[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a0a052b9 (
    .a(al_eb2ab31[21]),
    .b(al_8f688f54[21]),
    .c(al_ff6a88f6),
    .o({al_404f5287,al_e9628d6d[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b69c2ab8 (
    .a(al_eb2ab31[22]),
    .b(al_8f688f54[22]),
    .c(al_404f5287),
    .o({al_5d53cef6,al_e9628d6d[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_36356274 (
    .a(al_eb2ab31[23]),
    .b(al_8f688f54[23]),
    .c(al_5d53cef6),
    .o({al_4ed44021,al_e9628d6d[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d3d259de (
    .a(al_eb2ab31[24]),
    .b(al_8f688f54[24]),
    .c(al_4ed44021),
    .o({al_f392c8e6,al_e9628d6d[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_98c78a0d (
    .a(al_eb2ab31[25]),
    .b(al_8f688f54[25]),
    .c(al_f392c8e6),
    .o({al_cc8f42a5,al_e9628d6d[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2f204dfc (
    .a(al_eb2ab31[26]),
    .b(al_8f688f54[26]),
    .c(al_cc8f42a5),
    .o({al_3c97da5f,al_e9628d6d[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_83b3e627 (
    .a(al_eb2ab31[0]),
    .b(al_8f688f54[0]),
    .c(al_ca0ec285),
    .o({al_8a5edc6c,al_e9628d6d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2a2505ea (
    .a(al_eb2ab31[27]),
    .b(al_8f688f54[27]),
    .c(al_3c97da5f),
    .o({al_3bce7a34,al_e9628d6d[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a52b21c (
    .a(al_eb2ab31[28]),
    .b(al_8f688f54[28]),
    .c(al_3bce7a34),
    .o({open_n11,al_e9628d6d[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c85267b2 (
    .a(al_eb2ab31[1]),
    .b(al_8f688f54[1]),
    .c(al_8a5edc6c),
    .o({al_82b795a6,al_e9628d6d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2c6079d (
    .a(al_eb2ab31[2]),
    .b(al_8f688f54[2]),
    .c(al_82b795a6),
    .o({al_cb347ae8,al_e9628d6d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e5fbd1e5 (
    .a(al_eb2ab31[3]),
    .b(al_8f688f54[3]),
    .c(al_cb347ae8),
    .o({al_fbe9b8eb,al_e9628d6d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fe459258 (
    .a(al_eb2ab31[4]),
    .b(al_8f688f54[4]),
    .c(al_fbe9b8eb),
    .o({al_855a8144,al_e9628d6d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3492dd27 (
    .a(al_eb2ab31[5]),
    .b(al_8f688f54[5]),
    .c(al_855a8144),
    .o({al_50dcf253,al_e9628d6d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fb8b8bd8 (
    .a(al_eb2ab31[6]),
    .b(al_8f688f54[6]),
    .c(al_50dcf253),
    .o({al_5a7c92db,al_e9628d6d[6]}));
  AL_DFF_X al_7ead5a66 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[0]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[0]));
  AL_DFF_X al_af2172e3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[9]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[9]));
  AL_DFF_X al_c2e3ceaf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[10]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[10]));
  AL_DFF_X al_dc335f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[11]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[11]));
  AL_DFF_X al_ddeee205 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[12]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[12]));
  AL_DFF_X al_a19273e5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[13]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[13]));
  AL_DFF_X al_154ed596 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[14]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[14]));
  AL_DFF_X al_164c13ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[15]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[15]));
  AL_DFF_X al_e6352f12 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[16]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[16]));
  AL_DFF_X al_f5c5cb6b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[17]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[17]));
  AL_DFF_X al_ebc56e22 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[18]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[18]));
  AL_DFF_X al_e92df8f7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[1]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[1]));
  AL_DFF_X al_3c2569fd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[19]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[19]));
  AL_DFF_X al_7a198bed (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[20]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[20]));
  AL_DFF_X al_b227226b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[21]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[21]));
  AL_DFF_X al_6bb79861 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[22]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[22]));
  AL_DFF_X al_d8782f24 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[23]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[23]));
  AL_DFF_X al_e2551fd6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[24]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[24]));
  AL_DFF_X al_1404544f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[25]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[25]));
  AL_DFF_X al_c64ff9b3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[26]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[26]));
  AL_DFF_X al_4535f59d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[27]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[27]));
  AL_DFF_X al_83c74193 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[28]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[28]));
  AL_DFF_X al_cecc45f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[2]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[2]));
  AL_DFF_X al_2e824c2c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[3]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[3]));
  AL_DFF_X al_1cf54db9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[4]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[4]));
  AL_DFF_X al_f01e204a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[5]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[5]));
  AL_DFF_X al_24069c01 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[6]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[6]));
  AL_DFF_X al_4844f678 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[7]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[7]));
  AL_DFF_X al_5638f66b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_480f15b7[8]),
    .en(din_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eb2ab31[8]));
  AL_DFF_X al_ae00e8bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_54f6d4d2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_418f7602));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8cbdec3a (
    .a(al_8f688f54[7]),
    .b(al_4fe8581e[7]),
    .c(al_90fed4e7),
    .o({al_10238dc7,al_6d487ee0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2709750a (
    .a(al_8f688f54[8]),
    .b(al_4fe8581e[8]),
    .c(al_10238dc7),
    .o({al_8b4171c8,al_6d487ee0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_303f2f22 (
    .a(al_8f688f54[9]),
    .b(al_4fe8581e[9]),
    .c(al_8b4171c8),
    .o({al_2c346a44,al_6d487ee0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ef85db2d (
    .a(al_8f688f54[10]),
    .b(al_4fe8581e[10]),
    .c(al_2c346a44),
    .o({al_36624d30,al_6d487ee0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3c069ca7 (
    .a(al_8f688f54[11]),
    .b(al_4fe8581e[11]),
    .c(al_36624d30),
    .o({al_438b278b,al_6d487ee0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cb5efe90 (
    .a(al_8f688f54[12]),
    .b(al_4fe8581e[12]),
    .c(al_438b278b),
    .o({al_de0bda5,al_6d487ee0[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_727c48ae (
    .a(al_8f688f54[13]),
    .b(al_4fe8581e[13]),
    .c(al_de0bda5),
    .o({al_89db50f8,al_6d487ee0[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_90267592 (
    .a(al_8f688f54[14]),
    .b(al_4fe8581e[14]),
    .c(al_89db50f8),
    .o({al_d2835c11,al_6d487ee0[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_29dffe8d (
    .a(al_8f688f54[15]),
    .b(al_4fe8581e[15]),
    .c(al_d2835c11),
    .o({al_e0e4e676,al_6d487ee0[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_47f0b456 (
    .a(al_8f688f54[16]),
    .b(al_4fe8581e[16]),
    .c(al_e0e4e676),
    .o({al_685ac330,al_6d487ee0[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_790906ba (
    .a(1'b0),
    .o({al_dd04a5ca,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6023f309 (
    .a(al_8f688f54[17]),
    .b(al_4fe8581e[17]),
    .c(al_685ac330),
    .o({al_bc1a95db,al_6d487ee0[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4a423d0e (
    .a(al_8f688f54[18]),
    .b(al_4fe8581e[18]),
    .c(al_bc1a95db),
    .o({al_c7938c90,al_6d487ee0[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fbb5b95a (
    .a(al_8f688f54[19]),
    .b(al_4fe8581e[19]),
    .c(al_c7938c90),
    .o({al_3b1bd3d,al_6d487ee0[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_eb339349 (
    .a(al_8f688f54[20]),
    .b(al_4fe8581e[20]),
    .c(al_3b1bd3d),
    .o({al_1c7d78dc,al_6d487ee0[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dc0a517e (
    .a(al_8f688f54[21]),
    .b(al_4fe8581e[21]),
    .c(al_1c7d78dc),
    .o({al_c4c4b744,al_6d487ee0[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a63b0d7 (
    .a(al_8f688f54[22]),
    .b(al_4fe8581e[22]),
    .c(al_c4c4b744),
    .o({al_82fc816d,al_6d487ee0[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9b0f4d17 (
    .a(al_8f688f54[23]),
    .b(al_4fe8581e[23]),
    .c(al_82fc816d),
    .o({al_85782b8c,al_6d487ee0[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_afe55e8f (
    .a(al_8f688f54[24]),
    .b(al_4fe8581e[24]),
    .c(al_85782b8c),
    .o({al_52d5f2ec,al_6d487ee0[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1c952176 (
    .a(al_8f688f54[25]),
    .b(al_4fe8581e[25]),
    .c(al_52d5f2ec),
    .o({al_ce46c960,al_6d487ee0[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3e5f5426 (
    .a(al_8f688f54[26]),
    .b(al_4fe8581e[26]),
    .c(al_ce46c960),
    .o({al_8d67c17b,al_6d487ee0[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_370a3ed4 (
    .a(al_8f688f54[0]),
    .b(al_4fe8581e[0]),
    .c(al_dd04a5ca),
    .o({al_461ca1b0,al_6d487ee0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1265508c (
    .a(al_8f688f54[27]),
    .b(al_4fe8581e[27]),
    .c(al_8d67c17b),
    .o({al_6b121a3b,al_6d487ee0[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_beae7fc1 (
    .a(al_8f688f54[28]),
    .b(al_4fe8581e[28]),
    .c(al_6b121a3b),
    .o({open_n15,al_6d487ee0[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_80dc6f42 (
    .a(al_8f688f54[1]),
    .b(al_4fe8581e[1]),
    .c(al_461ca1b0),
    .o({al_dec8e5a2,al_6d487ee0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cbd79a66 (
    .a(al_8f688f54[2]),
    .b(al_4fe8581e[2]),
    .c(al_dec8e5a2),
    .o({al_66eadc2c,al_6d487ee0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_34d27e90 (
    .a(al_8f688f54[3]),
    .b(al_4fe8581e[3]),
    .c(al_66eadc2c),
    .o({al_60c7c36e,al_6d487ee0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b3b886c1 (
    .a(al_8f688f54[4]),
    .b(al_4fe8581e[4]),
    .c(al_60c7c36e),
    .o({al_8f3aa2df,al_6d487ee0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b17057c4 (
    .a(al_8f688f54[5]),
    .b(al_4fe8581e[5]),
    .c(al_8f3aa2df),
    .o({al_fb131175,al_6d487ee0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2696884a (
    .a(al_8f688f54[6]),
    .b(al_4fe8581e[6]),
    .c(al_fb131175),
    .o({al_90fed4e7,al_6d487ee0[6]}));
  AL_DFF_X al_11e34ed7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[0]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[0]));
  AL_DFF_X al_283840c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[9]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[9]));
  AL_DFF_X al_a9b8ce30 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[10]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[10]));
  AL_DFF_X al_df3578f2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[11]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[11]));
  AL_DFF_X al_a575c43a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[12]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[12]));
  AL_DFF_X al_2797f704 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[13]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[13]));
  AL_DFF_X al_b28bc32 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[14]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[14]));
  AL_DFF_X al_2ad57e11 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[15]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[15]));
  AL_DFF_X al_85624d35 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[16]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[16]));
  AL_DFF_X al_6132b32f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[17]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[17]));
  AL_DFF_X al_741ad1b7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[18]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[18]));
  AL_DFF_X al_f5b54ee6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[1]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[1]));
  AL_DFF_X al_cccedf51 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[19]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[19]));
  AL_DFF_X al_cd746bec (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[20]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[20]));
  AL_DFF_X al_bbbd528 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[21]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[21]));
  AL_DFF_X al_1cbf35e9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[22]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[22]));
  AL_DFF_X al_69415f6c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[23]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[23]));
  AL_DFF_X al_e3150e0e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[24]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[24]));
  AL_DFF_X al_98b9980e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[25]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[25]));
  AL_DFF_X al_1bf2d452 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[26]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[26]));
  AL_DFF_X al_abb73263 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[27]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[27]));
  AL_DFF_X al_87b4502d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[28]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[28]));
  AL_DFF_X al_264a2f27 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[2]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[2]));
  AL_DFF_X al_b021a5d0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[3]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[3]));
  AL_DFF_X al_38570098 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[4]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[4]));
  AL_DFF_X al_b95de5f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[5]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[5]));
  AL_DFF_X al_3413944a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[6]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[6]));
  AL_DFF_X al_3b9e7285 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[7]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[7]));
  AL_DFF_X al_18236158 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_e9628d6d[8]),
    .en(al_54f6d4d2),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f688f54[8]));
  AL_DFF_X al_b5b5360 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_418f7602),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2867582b));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_419a1774 (
    .a(al_4fe8581e[7]),
    .b(al_7d3eb7bc[7]),
    .c(al_31957fb7),
    .o({al_40f92736,al_feb3b069[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b695b53b (
    .a(al_4fe8581e[8]),
    .b(al_7d3eb7bc[8]),
    .c(al_40f92736),
    .o({al_bc0758d,al_feb3b069[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_db79f0c4 (
    .a(al_4fe8581e[9]),
    .b(al_7d3eb7bc[9]),
    .c(al_bc0758d),
    .o({al_98711f8a,al_feb3b069[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7456b95c (
    .a(al_4fe8581e[10]),
    .b(al_7d3eb7bc[10]),
    .c(al_98711f8a),
    .o({al_62e158f1,al_feb3b069[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_81a933c2 (
    .a(al_4fe8581e[11]),
    .b(al_7d3eb7bc[11]),
    .c(al_62e158f1),
    .o({al_bd8fc407,al_feb3b069[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_aa151bcb (
    .a(al_4fe8581e[12]),
    .b(al_7d3eb7bc[12]),
    .c(al_bd8fc407),
    .o({al_b1815462,al_feb3b069[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ab36186b (
    .a(al_4fe8581e[13]),
    .b(al_7d3eb7bc[13]),
    .c(al_b1815462),
    .o({al_e23d25b3,al_feb3b069[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9e805954 (
    .a(al_4fe8581e[14]),
    .b(al_7d3eb7bc[14]),
    .c(al_e23d25b3),
    .o({al_62be7f6f,al_feb3b069[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b7404e88 (
    .a(al_4fe8581e[15]),
    .b(al_7d3eb7bc[15]),
    .c(al_62be7f6f),
    .o({al_58af7ea5,al_feb3b069[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f3f9a8ab (
    .a(al_4fe8581e[16]),
    .b(al_7d3eb7bc[16]),
    .c(al_58af7ea5),
    .o({al_6b633f05,al_feb3b069[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_627b4658 (
    .a(1'b0),
    .o({al_62124ca0,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_404f0ebb (
    .a(al_4fe8581e[17]),
    .b(al_7d3eb7bc[17]),
    .c(al_6b633f05),
    .o({al_fcebab7e,al_feb3b069[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2b7458bb (
    .a(al_4fe8581e[18]),
    .b(al_7d3eb7bc[18]),
    .c(al_fcebab7e),
    .o({al_53c60bff,al_feb3b069[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f77f52cc (
    .a(al_4fe8581e[19]),
    .b(al_7d3eb7bc[19]),
    .c(al_53c60bff),
    .o({al_1b2cf291,al_feb3b069[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_80f5581d (
    .a(al_4fe8581e[20]),
    .b(al_7d3eb7bc[20]),
    .c(al_1b2cf291),
    .o({al_e060e572,al_feb3b069[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e92be987 (
    .a(al_4fe8581e[21]),
    .b(al_7d3eb7bc[21]),
    .c(al_e060e572),
    .o({al_d57ca002,al_feb3b069[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_201eb23f (
    .a(al_4fe8581e[22]),
    .b(al_7d3eb7bc[22]),
    .c(al_d57ca002),
    .o({al_9f2e787e,al_feb3b069[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a5a4b6ab (
    .a(al_4fe8581e[23]),
    .b(al_7d3eb7bc[23]),
    .c(al_9f2e787e),
    .o({al_560a769,al_feb3b069[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7b464882 (
    .a(al_4fe8581e[24]),
    .b(al_7d3eb7bc[24]),
    .c(al_560a769),
    .o({al_f76ae046,al_feb3b069[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a468c488 (
    .a(al_4fe8581e[25]),
    .b(al_7d3eb7bc[25]),
    .c(al_f76ae046),
    .o({al_1b884b48,al_feb3b069[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bcc58b03 (
    .a(al_4fe8581e[26]),
    .b(al_7d3eb7bc[26]),
    .c(al_1b884b48),
    .o({al_45855c0b,al_feb3b069[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d5ae9b55 (
    .a(al_4fe8581e[0]),
    .b(al_7d3eb7bc[0]),
    .c(al_62124ca0),
    .o({al_2e19f2fe,al_feb3b069[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_19452c6 (
    .a(al_4fe8581e[27]),
    .b(al_7d3eb7bc[27]),
    .c(al_45855c0b),
    .o({al_3a284b58,al_feb3b069[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_81f55882 (
    .a(al_4fe8581e[28]),
    .b(al_7d3eb7bc[28]),
    .c(al_3a284b58),
    .o({open_n19,al_feb3b069[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c5b727e7 (
    .a(al_4fe8581e[1]),
    .b(al_7d3eb7bc[1]),
    .c(al_2e19f2fe),
    .o({al_a1734311,al_feb3b069[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7c325c16 (
    .a(al_4fe8581e[2]),
    .b(al_7d3eb7bc[2]),
    .c(al_a1734311),
    .o({al_9b8ea422,al_feb3b069[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6f096261 (
    .a(al_4fe8581e[3]),
    .b(al_7d3eb7bc[3]),
    .c(al_9b8ea422),
    .o({al_d548edf7,al_feb3b069[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cc0b6c89 (
    .a(al_4fe8581e[4]),
    .b(al_7d3eb7bc[4]),
    .c(al_d548edf7),
    .o({al_6bb3744a,al_feb3b069[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_37dff7a1 (
    .a(al_4fe8581e[5]),
    .b(al_7d3eb7bc[5]),
    .c(al_6bb3744a),
    .o({al_70d5777e,al_feb3b069[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ca06cb4a (
    .a(al_4fe8581e[6]),
    .b(al_7d3eb7bc[6]),
    .c(al_70d5777e),
    .o({al_31957fb7,al_feb3b069[6]}));
  AL_DFF_X al_e11570b7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[0]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[0]));
  AL_DFF_X al_1d0efb82 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[9]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[9]));
  AL_DFF_X al_180d17 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[10]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[10]));
  AL_DFF_X al_73f17f4c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[11]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[11]));
  AL_DFF_X al_45dcf38f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[12]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[12]));
  AL_DFF_X al_29358c14 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[13]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[13]));
  AL_DFF_X al_168d471d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[14]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[14]));
  AL_DFF_X al_4e41950d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[15]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[15]));
  AL_DFF_X al_e1ed56ce (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[16]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[16]));
  AL_DFF_X al_b2ca9648 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[17]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[17]));
  AL_DFF_X al_69e6acab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[18]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[18]));
  AL_DFF_X al_96fb6dc6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[1]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[1]));
  AL_DFF_X al_73a06250 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[19]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[19]));
  AL_DFF_X al_e32b7ccc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[20]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[20]));
  AL_DFF_X al_2bfc91d8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[21]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[21]));
  AL_DFF_X al_b328303b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[22]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[22]));
  AL_DFF_X al_391ef9cc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[23]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[23]));
  AL_DFF_X al_5433ff1f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[24]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[24]));
  AL_DFF_X al_7715632a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[25]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[25]));
  AL_DFF_X al_35663785 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[26]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[26]));
  AL_DFF_X al_c39a6666 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[27]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[27]));
  AL_DFF_X al_e8ff3d24 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[28]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[28]));
  AL_DFF_X al_72ae767c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[2]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[2]));
  AL_DFF_X al_4effa87e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[3]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[3]));
  AL_DFF_X al_29ff22fa (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[4]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[4]));
  AL_DFF_X al_31402a33 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[5]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[5]));
  AL_DFF_X al_7cb6afde (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[6]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[6]));
  AL_DFF_X al_7b406089 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[7]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[7]));
  AL_DFF_X al_86762062 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_6d487ee0[8]),
    .en(al_418f7602),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fe8581e[8]));
  AL_DFF_X al_6b1c76f6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2867582b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b833a2e));
  AL_DFF_X al_2e35dc50 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[0]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[0]));
  AL_DFF_X al_b68b53b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[9]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[9]));
  AL_DFF_X al_b8ee8307 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[10]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[10]));
  AL_DFF_X al_f2d05973 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[11]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[11]));
  AL_DFF_X al_b3cf66d4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[12]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[12]));
  AL_DFF_X al_185e10fc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[13]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[13]));
  AL_DFF_X al_8b32e91f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[14]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[14]));
  AL_DFF_X al_1fa514ba (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[15]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[15]));
  AL_DFF_X al_78187ad9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[16]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[16]));
  AL_DFF_X al_a1a559a8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[17]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[17]));
  AL_DFF_X al_9afacfef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[18]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[18]));
  AL_DFF_X al_aad631cb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[1]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[1]));
  AL_DFF_X al_d44488ae (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[19]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[19]));
  AL_DFF_X al_8b2f80c1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[20]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[20]));
  AL_DFF_X al_e3674559 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[21]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[21]));
  AL_DFF_X al_c6ee3713 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[22]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[22]));
  AL_DFF_X al_5e078d4a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[23]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[23]));
  AL_DFF_X al_4320687d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[24]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[24]));
  AL_DFF_X al_3665567e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[25]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[25]));
  AL_DFF_X al_25aa00b8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[26]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[26]));
  AL_DFF_X al_e7e469af (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[27]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[27]));
  AL_DFF_X al_55f0b33c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[28]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[28]));
  AL_DFF_X al_865db970 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[2]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[2]));
  AL_DFF_X al_71e31c8e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[3]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[3]));
  AL_DFF_X al_d041ad2d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[4]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[4]));
  AL_DFF_X al_f52100be (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[5]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[5]));
  AL_DFF_X al_a12c0c0a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[6]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[6]));
  AL_DFF_X al_d05d0598 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[7]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[7]));
  AL_DFF_X al_b720a4a6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_feb3b069[8]),
    .en(al_2867582b),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d3eb7bc[8]));
  AL_DFF_X al_8a5c369b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[0]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[0]));
  AL_DFF_X al_e426e522 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[9]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[9]));
  AL_DFF_X al_88c76fb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[10]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[10]));
  AL_DFF_X al_5ee65d11 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[11]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[11]));
  AL_DFF_X al_930dd07d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[12]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[12]));
  AL_DFF_X al_8aabeb19 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[13]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[13]));
  AL_DFF_X al_d405111d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[14]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[14]));
  AL_DFF_X al_cd48a92e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[15]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[15]));
  AL_DFF_X al_5404bacc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[16]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[16]));
  AL_DFF_X al_a90e09b2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[17]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[17]));
  AL_DFF_X al_c0eb14a1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[18]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[18]));
  AL_DFF_X al_772b1557 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[1]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[1]));
  AL_DFF_X al_829c4174 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[19]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[19]));
  AL_DFF_X al_5e100677 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[20]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[20]));
  AL_DFF_X al_8fb1d0df (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[21]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[21]));
  AL_DFF_X al_57c89f56 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[22]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[22]));
  AL_DFF_X al_6b762143 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[23]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[23]));
  AL_DFF_X al_33d5049c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[24]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[24]));
  AL_DFF_X al_68d127bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[25]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[25]));
  AL_DFF_X al_b1a562ee (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[26]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[26]));
  AL_DFF_X al_987df877 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[27]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[27]));
  AL_DFF_X al_8d6b3342 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[28]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[28]));
  AL_DFF_X al_278bbfd4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[2]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[2]));
  AL_DFF_X al_37bddcac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[3]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[3]));
  AL_DFF_X al_49cfdb98 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[4]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[4]));
  AL_DFF_X al_21419022 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[5]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[5]));
  AL_DFF_X al_db7c9bef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[6]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[6]));
  AL_DFF_X al_d83b64ca (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[7]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[7]));
  AL_DFF_X al_82fbdbdb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c6636[8]),
    .en(al_8b833a2e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c916a43[8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_85829322 (
    .a(din_en),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .d(al_1deac949[2]),
    .o(al_65b98507));
  AL_DFF_X al_208ff28d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[0]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[0]));
  AL_DFF_X al_cb1a594d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[9]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[9]));
  AL_DFF_X al_59f2a9a0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[10]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[10]));
  AL_DFF_X al_84aec57d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[11]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[11]));
  AL_DFF_X al_6822c62f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[12]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[12]));
  AL_DFF_X al_ea7d814f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[13]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[13]));
  AL_DFF_X al_b98f781f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[14]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[14]));
  AL_DFF_X al_5ae5899a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[15]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[15]));
  AL_DFF_X al_9aa0a145 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[16]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[16]));
  AL_DFF_X al_fd6f5129 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[17]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[17]));
  AL_DFF_X al_8aca99a2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[18]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[18]));
  AL_DFF_X al_9cb79e4d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[1]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[1]));
  AL_DFF_X al_7686f558 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[19]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[19]));
  AL_DFF_X al_c5c1f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[20]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[20]));
  AL_DFF_X al_cc5d993d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[21]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[21]));
  AL_DFF_X al_13939656 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[22]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[22]));
  AL_DFF_X al_cdfdca31 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[23]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[23]));
  AL_DFF_X al_8ff91450 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[24]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[24]));
  AL_DFF_X al_975fc98b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[25]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[25]));
  AL_DFF_X al_dae2576b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[26]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[26]));
  AL_DFF_X al_a3e1a1e2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[27]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[27]));
  AL_DFF_X al_7e529903 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[28]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[28]));
  AL_DFF_X al_ccb7c64e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[2]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[2]));
  AL_DFF_X al_9c6b6b19 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[3]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[3]));
  AL_DFF_X al_95543770 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[4]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[4]));
  AL_DFF_X al_f8482182 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[5]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[5]));
  AL_DFF_X al_7d8e3654 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[6]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[6]));
  AL_DFF_X al_7d6ffb14 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[7]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[7]));
  AL_DFF_X al_c3fe3080 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2c916a43[8]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_62f4aab[8]));
  AL_DFF_X al_f4a7e0bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_65b98507),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3fe5f260));
  AL_DFF_X al_30fabc81 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[0]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[0]));
  AL_DFF_X al_9f453c00 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[9]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[9]));
  AL_DFF_X al_112d4d5a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[10]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[10]));
  AL_DFF_X al_97b196f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[11]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[11]));
  AL_DFF_X al_dbdd51a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[12]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[12]));
  AL_DFF_X al_ab193d58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[13]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[13]));
  AL_DFF_X al_3f89e8f3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[14]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[14]));
  AL_DFF_X al_75c709f7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[15]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[15]));
  AL_DFF_X al_92dbdb45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[16]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[16]));
  AL_DFF_X al_b083a1cd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[17]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[17]));
  AL_DFF_X al_2184ae49 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[18]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[18]));
  AL_DFF_X al_4f61e928 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[1]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[1]));
  AL_DFF_X al_b4eeed5e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[19]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[19]));
  AL_DFF_X al_a57f5a05 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[20]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[20]));
  AL_DFF_X al_daf88fa3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[21]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[21]));
  AL_DFF_X al_8c9cd5a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[22]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[22]));
  AL_DFF_X al_414d09fa (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[23]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[23]));
  AL_DFF_X al_9bf51a31 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[24]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[24]));
  AL_DFF_X al_e8777fdc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[25]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[25]));
  AL_DFF_X al_43f59c43 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[26]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[26]));
  AL_DFF_X al_e5c51b48 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[27]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[27]));
  AL_DFF_X al_d9bac04f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[28]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[28]));
  AL_DFF_X al_eee4ccbc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[2]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[2]));
  AL_DFF_X al_700234f3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[3]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[3]));
  AL_DFF_X al_3f290760 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[4]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[4]));
  AL_DFF_X al_3a8816a0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[5]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[5]));
  AL_DFF_X al_a4ad8988 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[6]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[6]));
  AL_DFF_X al_d5721ec9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[7]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[7]));
  AL_DFF_X al_47c13be9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4e1fa175[8]),
    .en(al_65b98507),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5414e669[8]));
  AL_DFF_X al_e8edcd6c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[0]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[0]));
  AL_DFF_X al_8918cf82 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[9]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[9]));
  AL_DFF_X al_1c612fa7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[10]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[10]));
  AL_DFF_X al_c21512c9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[11]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[11]));
  AL_DFF_X al_437f994c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[12]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[12]));
  AL_DFF_X al_63a15ae9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[13]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[13]));
  AL_DFF_X al_c2e857ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[14]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[14]));
  AL_DFF_X al_c87da315 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[15]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[15]));
  AL_DFF_X al_64619a0e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[16]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[16]));
  AL_DFF_X al_13ddf83c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[17]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[17]));
  AL_DFF_X al_ffec4da8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[18]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[18]));
  AL_DFF_X al_e58841b5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[1]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[1]));
  AL_DFF_X al_933707d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[19]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[19]));
  AL_DFF_X al_7e586ab4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[20]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[20]));
  AL_DFF_X al_f87d458c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[21]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[21]));
  AL_DFF_X al_56e8a919 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[22]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[22]));
  AL_DFF_X al_343113c8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[23]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[23]));
  AL_DFF_X al_e2268dc5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[24]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[24]));
  AL_DFF_X al_e6c50fdb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[25]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[25]));
  AL_DFF_X al_37f86324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[26]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[26]));
  AL_DFF_X al_28489c59 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[27]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[27]));
  AL_DFF_X al_23dbd431 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[28]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[28]));
  AL_DFF_X al_d244ccce (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[2]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[2]));
  AL_DFF_X al_cff09ca1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[3]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[3]));
  AL_DFF_X al_5a650fc7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[4]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[4]));
  AL_DFF_X al_bf1243d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[5]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[5]));
  AL_DFF_X al_f32b8273 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[6]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[6]));
  AL_DFF_X al_a522a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[7]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[7]));
  AL_DFF_X al_72325d94 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5414e669[8]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd893e44[8]));
  AL_DFF_X al_3e1a344a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3fe5f260),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81c141dd));
  AL_DFF_X al_7d302633 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[0]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[0]));
  AL_DFF_X al_3e889b8b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[9]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[9]));
  AL_DFF_X al_bb376bfe (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[10]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[10]));
  AL_DFF_X al_92fa971d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[11]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[11]));
  AL_DFF_X al_6050e582 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[12]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[12]));
  AL_DFF_X al_de6806a9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[13]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[13]));
  AL_DFF_X al_e979a902 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[14]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[14]));
  AL_DFF_X al_ecd4cd0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[15]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[15]));
  AL_DFF_X al_3265c949 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[16]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[16]));
  AL_DFF_X al_83a84588 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[17]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[17]));
  AL_DFF_X al_2d74a7c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[18]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[18]));
  AL_DFF_X al_fd07722d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[1]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[1]));
  AL_DFF_X al_5fec5d87 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[19]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[19]));
  AL_DFF_X al_1d813794 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[20]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[20]));
  AL_DFF_X al_abf61600 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[21]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[21]));
  AL_DFF_X al_8f441c6c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[22]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[22]));
  AL_DFF_X al_7d7562d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[23]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[23]));
  AL_DFF_X al_9ce52bbe (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[24]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[24]));
  AL_DFF_X al_c8e20e09 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[25]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[25]));
  AL_DFF_X al_e632b320 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[26]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[26]));
  AL_DFF_X al_912236d8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[27]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[27]));
  AL_DFF_X al_ac2d628e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[28]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[28]));
  AL_DFF_X al_49b1f36d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[2]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[2]));
  AL_DFF_X al_9cd8208f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[3]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[3]));
  AL_DFF_X al_89cbc291 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[4]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[4]));
  AL_DFF_X al_1094fdd3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[5]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[5]));
  AL_DFF_X al_483c3bcf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[6]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[6]));
  AL_DFF_X al_6da0d01 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[7]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[7]));
  AL_DFF_X al_51df0663 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4873fb93[8]),
    .en(al_3fe5f260),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b27b90b2[8]));
  AL_DFF_X al_e74b2f2a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[0]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[0]));
  AL_DFF_X al_75956fb7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[9]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[9]));
  AL_DFF_X al_86bc42e7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[10]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[10]));
  AL_DFF_X al_ab98a49b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[11]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[11]));
  AL_DFF_X al_d8ec79a1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[12]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[12]));
  AL_DFF_X al_59f3e5c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[13]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[13]));
  AL_DFF_X al_7f0a0d25 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[14]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[14]));
  AL_DFF_X al_600f72ea (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[15]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[15]));
  AL_DFF_X al_52030c86 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[16]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[16]));
  AL_DFF_X al_e4fccc3c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[17]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[17]));
  AL_DFF_X al_89b30cf8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[18]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[18]));
  AL_DFF_X al_b1fe82e2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[1]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[1]));
  AL_DFF_X al_a32b6b55 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[19]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[19]));
  AL_DFF_X al_44805624 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[20]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[20]));
  AL_DFF_X al_295838d0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[21]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[21]));
  AL_DFF_X al_fe1f4edf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[22]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[22]));
  AL_DFF_X al_23be9e97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[23]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[23]));
  AL_DFF_X al_3d0b697e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[24]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[24]));
  AL_DFF_X al_185b9fca (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[25]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[25]));
  AL_DFF_X al_b263a3f9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[26]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[26]));
  AL_DFF_X al_c12020b5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[27]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[27]));
  AL_DFF_X al_98118c1e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[28]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[28]));
  AL_DFF_X al_95a2c788 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[2]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[2]));
  AL_DFF_X al_fb3f37ad (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[3]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[3]));
  AL_DFF_X al_d4e2ca91 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[4]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[4]));
  AL_DFF_X al_9480b797 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[5]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[5]));
  AL_DFF_X al_48b506f7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[6]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[6]));
  AL_DFF_X al_178207c3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[7]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[7]));
  AL_DFF_X al_561a2de7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_b27b90b2[8]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9955f70[8]));
  AL_DFF_X al_ec2afc84 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_81c141dd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fd840f8c));
  AL_DFF_X al_27457f27 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[0]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[0]));
  AL_DFF_X al_df7e3663 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[9]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[9]));
  AL_DFF_X al_c005214 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[10]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[10]));
  AL_DFF_X al_50c33a4b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[11]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[11]));
  AL_DFF_X al_e36fc598 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[12]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[12]));
  AL_DFF_X al_42d8c3cc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[13]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[13]));
  AL_DFF_X al_748f74eb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[14]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[14]));
  AL_DFF_X al_bf58ea1f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[15]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[15]));
  AL_DFF_X al_89219365 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[16]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[16]));
  AL_DFF_X al_6420a58 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[17]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[17]));
  AL_DFF_X al_568a5e41 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[18]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[18]));
  AL_DFF_X al_49f9a2cd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[1]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[1]));
  AL_DFF_X al_c45a82ce (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[19]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[19]));
  AL_DFF_X al_ee81b4f0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[20]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[20]));
  AL_DFF_X al_d0fed496 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[21]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[21]));
  AL_DFF_X al_ce4f487d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[22]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[22]));
  AL_DFF_X al_f55c97e2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[23]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[23]));
  AL_DFF_X al_6d6b9d06 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[24]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[24]));
  AL_DFF_X al_1e129b6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[25]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[25]));
  AL_DFF_X al_d1517861 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[26]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[26]));
  AL_DFF_X al_edc2093f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[27]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[27]));
  AL_DFF_X al_9334945b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[28]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[28]));
  AL_DFF_X al_f667965c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[2]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[2]));
  AL_DFF_X al_bd3d00ba (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[3]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[3]));
  AL_DFF_X al_d6352aaa (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[4]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[4]));
  AL_DFF_X al_80a0e8e6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[5]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[5]));
  AL_DFF_X al_e8e50eb8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[6]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[6]));
  AL_DFF_X al_557f6a55 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[7]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[7]));
  AL_DFF_X al_59c3f030 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d9b93292[8]),
    .en(al_81c141dd),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14ec71c5[8]));
  AL_DFF_X al_734647a4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[0]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[0]));
  AL_DFF_X al_655568c0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[9]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[9]));
  AL_DFF_X al_85e5b876 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[10]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[10]));
  AL_DFF_X al_5bef718b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[11]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[11]));
  AL_DFF_X al_df27589f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[12]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[12]));
  AL_DFF_X al_b538b123 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[13]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[13]));
  AL_DFF_X al_b13bf8ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[14]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[14]));
  AL_DFF_X al_c219bab9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[15]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[15]));
  AL_DFF_X al_9ce16a35 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[16]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[16]));
  AL_DFF_X al_f1a8fcf3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[17]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[17]));
  AL_DFF_X al_1363329 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[18]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[18]));
  AL_DFF_X al_98d2e5fc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[1]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[1]));
  AL_DFF_X al_d1022d01 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[19]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[19]));
  AL_DFF_X al_f83457a3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[20]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[20]));
  AL_DFF_X al_ac4524ab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[21]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[21]));
  AL_DFF_X al_89ed1fb7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[22]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[22]));
  AL_DFF_X al_e09f5ff6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[23]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[23]));
  AL_DFF_X al_ad5bfcdf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[24]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[24]));
  AL_DFF_X al_ea3f22e9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[25]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[25]));
  AL_DFF_X al_83061b1c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[26]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[26]));
  AL_DFF_X al_c2c7e2f0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[27]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[27]));
  AL_DFF_X al_1b787f56 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[28]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[28]));
  AL_DFF_X al_e118d9a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[2]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[2]));
  AL_DFF_X al_b79c06b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[3]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[3]));
  AL_DFF_X al_cc4b3c54 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[4]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[4]));
  AL_DFF_X al_7289a038 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[5]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[5]));
  AL_DFF_X al_cd8fd1ae (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[6]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[6]));
  AL_DFF_X al_ad559718 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[7]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[7]));
  AL_DFF_X al_7f814cc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_14ec71c5[8]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_afdc4416[8]));
  AL_DFF_X al_b69436bd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_fd840f8c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4705248d));
  AL_DFF_X al_a133c6a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[0]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[0]));
  AL_DFF_X al_934991f5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[9]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[9]));
  AL_DFF_X al_bbb38589 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[10]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[10]));
  AL_DFF_X al_a7310234 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[11]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[11]));
  AL_DFF_X al_dc2f9380 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[12]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[12]));
  AL_DFF_X al_282d141 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[13]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[13]));
  AL_DFF_X al_87c4bc47 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[14]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[14]));
  AL_DFF_X al_3f7713da (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[15]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[15]));
  AL_DFF_X al_e8549816 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[16]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[16]));
  AL_DFF_X al_2b258fef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[17]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[17]));
  AL_DFF_X al_d03b1959 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[18]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[18]));
  AL_DFF_X al_2dfa4dd1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[1]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[1]));
  AL_DFF_X al_b47ba9c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[19]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[19]));
  AL_DFF_X al_185b092d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[20]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[20]));
  AL_DFF_X al_51b4b32b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[21]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[21]));
  AL_DFF_X al_5b6e4b16 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[22]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[22]));
  AL_DFF_X al_d771c413 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[23]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[23]));
  AL_DFF_X al_4c6c30a2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[24]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[24]));
  AL_DFF_X al_ba2c0379 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[25]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[25]));
  AL_DFF_X al_3fe74565 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[26]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[26]));
  AL_DFF_X al_6c3cd82b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[27]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[27]));
  AL_DFF_X al_e139ffab (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[28]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[28]));
  AL_DFF_X al_4f81bf48 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[2]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[2]));
  AL_DFF_X al_eabc5e55 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[3]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[3]));
  AL_DFF_X al_fea7d8eb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[4]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[4]));
  AL_DFF_X al_950b43d8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[5]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[5]));
  AL_DFF_X al_18e101d2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[6]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[6]));
  AL_DFF_X al_fe4b421c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[7]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[7]));
  AL_DFF_X al_a934d6c5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1d216208[8]),
    .en(al_fd840f8c),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e11d7be[8]));
  AL_DFF_X al_edd72b25 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[0]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[0]));
  AL_DFF_X al_73f81613 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[9]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[9]));
  AL_DFF_X al_1239143 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[10]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[10]));
  AL_DFF_X al_4cd3c09c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[11]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[11]));
  AL_DFF_X al_862cd9a0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[12]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[12]));
  AL_DFF_X al_a93f492c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[13]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[13]));
  AL_DFF_X al_cfb3897d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[14]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[14]));
  AL_DFF_X al_cbda9c7f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[15]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[15]));
  AL_DFF_X al_a4caa0a2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[16]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[16]));
  AL_DFF_X al_185950b6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[17]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[17]));
  AL_DFF_X al_35b537f4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[18]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[18]));
  AL_DFF_X al_75cbcebc (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[1]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[1]));
  AL_DFF_X al_91c17854 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[19]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[19]));
  AL_DFF_X al_c5ebfd2a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[20]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[20]));
  AL_DFF_X al_d854bcd2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[21]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[21]));
  AL_DFF_X al_69f4d2e9 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[22]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[22]));
  AL_DFF_X al_460ba6c1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[23]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[23]));
  AL_DFF_X al_c9e93a32 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[24]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[24]));
  AL_DFF_X al_43be7412 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[25]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[25]));
  AL_DFF_X al_2cc84a36 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[26]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[26]));
  AL_DFF_X al_d2fd6557 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[27]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[27]));
  AL_DFF_X al_531e5e72 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[28]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[28]));
  AL_DFF_X al_94a0c85b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[2]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[2]));
  AL_DFF_X al_cc37547a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[3]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[3]));
  AL_DFF_X al_d92047d3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[4]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[4]));
  AL_DFF_X al_cb2d2202 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[5]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[5]));
  AL_DFF_X al_c85c6be8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[6]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[6]));
  AL_DFF_X al_ef8dc198 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[7]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[7]));
  AL_DFF_X al_b3acc32e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_5e11d7be[8]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6d689829[8]));
  AL_DFF_X al_47b0ff5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_4705248d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_229e7e2c));
  AL_DFF_X al_1b81f7d5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[0]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[0]));
  AL_DFF_X al_cdaad52d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[9]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[9]));
  AL_DFF_X al_306c843a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[10]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[10]));
  AL_DFF_X al_c02d08f2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[11]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[11]));
  AL_DFF_X al_4bc4745a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[12]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[12]));
  AL_DFF_X al_75aa000e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[13]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[13]));
  AL_DFF_X al_70220b86 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[14]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[14]));
  AL_DFF_X al_58a7fec5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[15]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[15]));
  AL_DFF_X al_41534214 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[16]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[16]));
  AL_DFF_X al_888be32e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[17]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[17]));
  AL_DFF_X al_91a1abe2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[18]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[18]));
  AL_DFF_X al_86c112e4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[1]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[1]));
  AL_DFF_X al_dd722ad0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[19]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[19]));
  AL_DFF_X al_6c38572e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[20]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[20]));
  AL_DFF_X al_c50eef39 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[21]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[21]));
  AL_DFF_X al_631fdbb1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[22]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[22]));
  AL_DFF_X al_8d043f1d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[23]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[23]));
  AL_DFF_X al_8b71dede (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[24]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[24]));
  AL_DFF_X al_aa40f684 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[25]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[25]));
  AL_DFF_X al_c1ced9f1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[26]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[26]));
  AL_DFF_X al_4ec8fc67 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[27]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[27]));
  AL_DFF_X al_f724eb55 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[28]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[28]));
  AL_DFF_X al_a75532a5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[2]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[2]));
  AL_DFF_X al_4a6d3f23 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[3]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[3]));
  AL_DFF_X al_f66a0d66 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[4]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[4]));
  AL_DFF_X al_82e8dfec (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[5]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[5]));
  AL_DFF_X al_6bae4afe (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[6]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[6]));
  AL_DFF_X al_23ad83db (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[7]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[7]));
  AL_DFF_X al_4daf1426 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_ac1e65eb[8]),
    .en(al_4705248d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1358e4cb[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_3731118c (
    .a(1'b0),
    .o({al_ea32c6e1,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_5414e669[8]),
    .b(al_cd893e44[8]),
    .c(al_ca5b12bc),
    .o({al_b49c276a,al_4873fb93[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_5414e669[9]),
    .b(al_cd893e44[9]),
    .c(al_b49c276a),
    .o({al_a23af5a4,al_4873fb93[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_5414e669[10]),
    .b(al_cd893e44[10]),
    .c(al_a23af5a4),
    .o({al_fe2986b6,al_4873fb93[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_5414e669[11]),
    .b(al_cd893e44[11]),
    .c(al_fe2986b6),
    .o({al_875c79d9,al_4873fb93[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_5414e669[12]),
    .b(al_cd893e44[12]),
    .c(al_875c79d9),
    .o({al_d21ff3d4,al_4873fb93[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_5414e669[13]),
    .b(al_cd893e44[13]),
    .c(al_d21ff3d4),
    .o({al_20da7cd1,al_4873fb93[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_5414e669[14]),
    .b(al_cd893e44[14]),
    .c(al_20da7cd1),
    .o({al_4b6c2990,al_4873fb93[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_5414e669[15]),
    .b(al_cd893e44[15]),
    .c(al_4b6c2990),
    .o({al_2a9315a6,al_4873fb93[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_5414e669[16]),
    .b(al_cd893e44[16]),
    .c(al_2a9315a6),
    .o({al_b9c5d958,al_4873fb93[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_5414e669[17]),
    .b(al_cd893e44[17]),
    .c(al_b9c5d958),
    .o({al_56630a35,al_4873fb93[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5224f5b (
    .a(al_5414e669[0]),
    .b(al_cd893e44[0]),
    .c(al_ea32c6e1),
    .o({al_2ac97405,al_4873fb93[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_5414e669[18]),
    .b(al_cd893e44[18]),
    .c(al_56630a35),
    .o({al_a1b0b17a,al_4873fb93[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_5414e669[19]),
    .b(al_cd893e44[19]),
    .c(al_a1b0b17a),
    .o({al_7b07bb65,al_4873fb93[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_5414e669[20]),
    .b(al_cd893e44[20]),
    .c(al_7b07bb65),
    .o({al_9df2af8f,al_4873fb93[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_5414e669[21]),
    .b(al_cd893e44[21]),
    .c(al_9df2af8f),
    .o({al_df20ca5b,al_4873fb93[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_5414e669[22]),
    .b(al_cd893e44[22]),
    .c(al_df20ca5b),
    .o({al_ab6a0e7,al_4873fb93[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e359bb16 (
    .a(al_5414e669[23]),
    .b(al_cd893e44[23]),
    .c(al_ab6a0e7),
    .o({al_3f047599,al_4873fb93[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6af83b3 (
    .a(al_5414e669[24]),
    .b(al_cd893e44[24]),
    .c(al_3f047599),
    .o({al_b4d1b2a2,al_4873fb93[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_717da7cc (
    .a(al_5414e669[25]),
    .b(al_cd893e44[25]),
    .c(al_b4d1b2a2),
    .o({al_469cb985,al_4873fb93[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_916a9569 (
    .a(al_5414e669[26]),
    .b(al_cd893e44[26]),
    .c(al_469cb985),
    .o({al_ffb568cb,al_4873fb93[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b53f57fa (
    .a(al_5414e669[27]),
    .b(al_cd893e44[27]),
    .c(al_ffb568cb),
    .o({al_8f0bd67f,al_4873fb93[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_5414e669[1]),
    .b(al_cd893e44[1]),
    .c(al_2ac97405),
    .o({al_a0ebd25,al_4873fb93[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_edf2dc1f (
    .a(al_5414e669[28]),
    .b(al_cd893e44[28]),
    .c(al_8f0bd67f),
    .o({open_n23,al_4873fb93[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_5414e669[2]),
    .b(al_cd893e44[2]),
    .c(al_a0ebd25),
    .o({al_f77a35ee,al_4873fb93[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_5414e669[3]),
    .b(al_cd893e44[3]),
    .c(al_f77a35ee),
    .o({al_2902a00c,al_4873fb93[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_5414e669[4]),
    .b(al_cd893e44[4]),
    .c(al_2902a00c),
    .o({al_94925fa9,al_4873fb93[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_5414e669[5]),
    .b(al_cd893e44[5]),
    .c(al_94925fa9),
    .o({al_51a70210,al_4873fb93[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_5414e669[6]),
    .b(al_cd893e44[6]),
    .c(al_51a70210),
    .o({al_fbeca432,al_4873fb93[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_5414e669[7]),
    .b(al_cd893e44[7]),
    .c(al_fbeca432),
    .o({al_ca5b12bc,al_4873fb93[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_3a3a68e0 (
    .a(1'b0),
    .o({al_b0d09b8,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7a9fe52 (
    .a(al_b27b90b2[8]),
    .b(al_9955f70[8]),
    .c(al_1e9cae1d),
    .o({al_13006735,al_d9b93292[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5542edfe (
    .a(al_b27b90b2[9]),
    .b(al_9955f70[9]),
    .c(al_13006735),
    .o({al_bbd9355,al_d9b93292[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_488602ff (
    .a(al_b27b90b2[10]),
    .b(al_9955f70[10]),
    .c(al_bbd9355),
    .o({al_8f481ef9,al_d9b93292[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e1d0a51 (
    .a(al_b27b90b2[11]),
    .b(al_9955f70[11]),
    .c(al_8f481ef9),
    .o({al_9ab66270,al_d9b93292[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a28406e8 (
    .a(al_b27b90b2[12]),
    .b(al_9955f70[12]),
    .c(al_9ab66270),
    .o({al_4dcb26fa,al_d9b93292[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b74b0b2 (
    .a(al_b27b90b2[13]),
    .b(al_9955f70[13]),
    .c(al_4dcb26fa),
    .o({al_d0181d13,al_d9b93292[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_225d9869 (
    .a(al_b27b90b2[14]),
    .b(al_9955f70[14]),
    .c(al_d0181d13),
    .o({al_b08aad73,al_d9b93292[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57140763 (
    .a(al_b27b90b2[15]),
    .b(al_9955f70[15]),
    .c(al_b08aad73),
    .o({al_c1c08587,al_d9b93292[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2faa1616 (
    .a(al_b27b90b2[16]),
    .b(al_9955f70[16]),
    .c(al_c1c08587),
    .o({al_689cec14,al_d9b93292[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed62317d (
    .a(al_b27b90b2[17]),
    .b(al_9955f70[17]),
    .c(al_689cec14),
    .o({al_9ddddc8e,al_d9b93292[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5194f578 (
    .a(al_b27b90b2[0]),
    .b(al_9955f70[0]),
    .c(al_b0d09b8),
    .o({al_94c23594,al_d9b93292[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd47866c (
    .a(al_b27b90b2[18]),
    .b(al_9955f70[18]),
    .c(al_9ddddc8e),
    .o({al_41a92fc7,al_d9b93292[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de077e95 (
    .a(al_b27b90b2[19]),
    .b(al_9955f70[19]),
    .c(al_41a92fc7),
    .o({al_d4d70e4b,al_d9b93292[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ff0b0f0 (
    .a(al_b27b90b2[20]),
    .b(al_9955f70[20]),
    .c(al_d4d70e4b),
    .o({al_e800c9ef,al_d9b93292[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84a7f2c5 (
    .a(al_b27b90b2[21]),
    .b(al_9955f70[21]),
    .c(al_e800c9ef),
    .o({al_5cf39772,al_d9b93292[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd22e386 (
    .a(al_b27b90b2[22]),
    .b(al_9955f70[22]),
    .c(al_5cf39772),
    .o({al_339b3bc,al_d9b93292[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e9daf8ce (
    .a(al_b27b90b2[23]),
    .b(al_9955f70[23]),
    .c(al_339b3bc),
    .o({al_c6da537,al_d9b93292[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b718cdc3 (
    .a(al_b27b90b2[24]),
    .b(al_9955f70[24]),
    .c(al_c6da537),
    .o({al_35361f12,al_d9b93292[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_220d3472 (
    .a(al_b27b90b2[25]),
    .b(al_9955f70[25]),
    .c(al_35361f12),
    .o({al_c6028b1e,al_d9b93292[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_446777ef (
    .a(al_b27b90b2[26]),
    .b(al_9955f70[26]),
    .c(al_c6028b1e),
    .o({al_87b345e3,al_d9b93292[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a586468 (
    .a(al_b27b90b2[27]),
    .b(al_9955f70[27]),
    .c(al_87b345e3),
    .o({al_29505f4f,al_d9b93292[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5250c82 (
    .a(al_b27b90b2[1]),
    .b(al_9955f70[1]),
    .c(al_94c23594),
    .o({al_d203b819,al_d9b93292[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e9578c63 (
    .a(al_b27b90b2[28]),
    .b(al_9955f70[28]),
    .c(al_29505f4f),
    .o({open_n27,al_d9b93292[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce5b7c47 (
    .a(al_b27b90b2[2]),
    .b(al_9955f70[2]),
    .c(al_d203b819),
    .o({al_c5f97e65,al_d9b93292[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2348e63f (
    .a(al_b27b90b2[3]),
    .b(al_9955f70[3]),
    .c(al_c5f97e65),
    .o({al_5aa7ca6a,al_d9b93292[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1dde6515 (
    .a(al_b27b90b2[4]),
    .b(al_9955f70[4]),
    .c(al_5aa7ca6a),
    .o({al_c709f85a,al_d9b93292[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_730170d3 (
    .a(al_b27b90b2[5]),
    .b(al_9955f70[5]),
    .c(al_c709f85a),
    .o({al_26a0aae,al_d9b93292[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_81729e9d (
    .a(al_b27b90b2[6]),
    .b(al_9955f70[6]),
    .c(al_26a0aae),
    .o({al_94b1300d,al_d9b93292[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73503454 (
    .a(al_b27b90b2[7]),
    .b(al_9955f70[7]),
    .c(al_94b1300d),
    .o({al_1e9cae1d,al_d9b93292[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_69abf9ec (
    .a(1'b0),
    .o({al_aa8f2cd8,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dfdc771 (
    .a(al_14ec71c5[8]),
    .b(al_afdc4416[8]),
    .c(al_16b99b31),
    .o({al_5c3c8bc3,al_1d216208[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e93dcd8b (
    .a(al_14ec71c5[9]),
    .b(al_afdc4416[9]),
    .c(al_5c3c8bc3),
    .o({al_83d3841d,al_1d216208[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f94769 (
    .a(al_14ec71c5[10]),
    .b(al_afdc4416[10]),
    .c(al_83d3841d),
    .o({al_21712447,al_1d216208[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18f640ef (
    .a(al_14ec71c5[11]),
    .b(al_afdc4416[11]),
    .c(al_21712447),
    .o({al_e26baa7c,al_1d216208[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86ec8670 (
    .a(al_14ec71c5[12]),
    .b(al_afdc4416[12]),
    .c(al_e26baa7c),
    .o({al_bd632267,al_1d216208[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6df03772 (
    .a(al_14ec71c5[13]),
    .b(al_afdc4416[13]),
    .c(al_bd632267),
    .o({al_7b0a2fb3,al_1d216208[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45f02cda (
    .a(al_14ec71c5[14]),
    .b(al_afdc4416[14]),
    .c(al_7b0a2fb3),
    .o({al_b8ace6d9,al_1d216208[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6b2c7c5 (
    .a(al_14ec71c5[15]),
    .b(al_afdc4416[15]),
    .c(al_b8ace6d9),
    .o({al_18580a3b,al_1d216208[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f06d29 (
    .a(al_14ec71c5[16]),
    .b(al_afdc4416[16]),
    .c(al_18580a3b),
    .o({al_830367be,al_1d216208[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff64c9f9 (
    .a(al_14ec71c5[17]),
    .b(al_afdc4416[17]),
    .c(al_830367be),
    .o({al_92e30c9d,al_1d216208[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6219435f (
    .a(al_14ec71c5[0]),
    .b(al_afdc4416[0]),
    .c(al_aa8f2cd8),
    .o({al_685d248f,al_1d216208[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_689e06a4 (
    .a(al_14ec71c5[18]),
    .b(al_afdc4416[18]),
    .c(al_92e30c9d),
    .o({al_6566c57e,al_1d216208[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a011db00 (
    .a(al_14ec71c5[19]),
    .b(al_afdc4416[19]),
    .c(al_6566c57e),
    .o({al_29ad0e3a,al_1d216208[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebcca0b3 (
    .a(al_14ec71c5[20]),
    .b(al_afdc4416[20]),
    .c(al_29ad0e3a),
    .o({al_51513f80,al_1d216208[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b00f8a2c (
    .a(al_14ec71c5[21]),
    .b(al_afdc4416[21]),
    .c(al_51513f80),
    .o({al_1cd5a819,al_1d216208[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67573096 (
    .a(al_14ec71c5[22]),
    .b(al_afdc4416[22]),
    .c(al_1cd5a819),
    .o({al_11e537d,al_1d216208[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a4bf0f3d (
    .a(al_14ec71c5[23]),
    .b(al_afdc4416[23]),
    .c(al_11e537d),
    .o({al_5d5b70cd,al_1d216208[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4075baa3 (
    .a(al_14ec71c5[24]),
    .b(al_afdc4416[24]),
    .c(al_5d5b70cd),
    .o({al_397e2eb4,al_1d216208[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68c3dc57 (
    .a(al_14ec71c5[25]),
    .b(al_afdc4416[25]),
    .c(al_397e2eb4),
    .o({al_60062243,al_1d216208[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac251091 (
    .a(al_14ec71c5[26]),
    .b(al_afdc4416[26]),
    .c(al_60062243),
    .o({al_14a9163b,al_1d216208[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f80b960 (
    .a(al_14ec71c5[27]),
    .b(al_afdc4416[27]),
    .c(al_14a9163b),
    .o({al_ca0bd035,al_1d216208[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9173b3c2 (
    .a(al_14ec71c5[1]),
    .b(al_afdc4416[1]),
    .c(al_685d248f),
    .o({al_cfde68ec,al_1d216208[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_798abbb4 (
    .a(al_14ec71c5[28]),
    .b(al_afdc4416[28]),
    .c(al_ca0bd035),
    .o({open_n31,al_1d216208[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e14f1c1 (
    .a(al_14ec71c5[2]),
    .b(al_afdc4416[2]),
    .c(al_cfde68ec),
    .o({al_5c1d9288,al_1d216208[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b174dbc (
    .a(al_14ec71c5[3]),
    .b(al_afdc4416[3]),
    .c(al_5c1d9288),
    .o({al_1f7974b0,al_1d216208[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6657a45b (
    .a(al_14ec71c5[4]),
    .b(al_afdc4416[4]),
    .c(al_1f7974b0),
    .o({al_c964d6b6,al_1d216208[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17e08140 (
    .a(al_14ec71c5[5]),
    .b(al_afdc4416[5]),
    .c(al_c964d6b6),
    .o({al_d5344387,al_1d216208[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e94e10ff (
    .a(al_14ec71c5[6]),
    .b(al_afdc4416[6]),
    .c(al_d5344387),
    .o({al_944a7435,al_1d216208[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_440a3abe (
    .a(al_14ec71c5[7]),
    .b(al_afdc4416[7]),
    .c(al_944a7435),
    .o({al_16b99b31,al_1d216208[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1e5edfe5 (
    .a(1'b0),
    .o({al_10ad2d4,open_n34}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d97c2b0d (
    .a(al_5e11d7be[8]),
    .b(al_6d689829[8]),
    .c(al_74c02a6e),
    .o({al_2c19a30d,al_ac1e65eb[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b7d12a4 (
    .a(al_5e11d7be[9]),
    .b(al_6d689829[9]),
    .c(al_2c19a30d),
    .o({al_30e98b36,al_ac1e65eb[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fb59cdb6 (
    .a(al_5e11d7be[10]),
    .b(al_6d689829[10]),
    .c(al_30e98b36),
    .o({al_dff2b81e,al_ac1e65eb[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_366a9dbb (
    .a(al_5e11d7be[11]),
    .b(al_6d689829[11]),
    .c(al_dff2b81e),
    .o({al_7e683184,al_ac1e65eb[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4a192c65 (
    .a(al_5e11d7be[12]),
    .b(al_6d689829[12]),
    .c(al_7e683184),
    .o({al_b5ad59ae,al_ac1e65eb[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_264762b0 (
    .a(al_5e11d7be[13]),
    .b(al_6d689829[13]),
    .c(al_b5ad59ae),
    .o({al_fdc784df,al_ac1e65eb[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a245e86f (
    .a(al_5e11d7be[14]),
    .b(al_6d689829[14]),
    .c(al_fdc784df),
    .o({al_8625eee6,al_ac1e65eb[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_361c4f76 (
    .a(al_5e11d7be[15]),
    .b(al_6d689829[15]),
    .c(al_8625eee6),
    .o({al_b46339ca,al_ac1e65eb[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_76a00777 (
    .a(al_5e11d7be[16]),
    .b(al_6d689829[16]),
    .c(al_b46339ca),
    .o({al_47553d9c,al_ac1e65eb[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fb02f698 (
    .a(al_5e11d7be[17]),
    .b(al_6d689829[17]),
    .c(al_47553d9c),
    .o({al_e55eeb92,al_ac1e65eb[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_28abd0a1 (
    .a(al_5e11d7be[0]),
    .b(al_6d689829[0]),
    .c(al_10ad2d4),
    .o({al_4b7e6f4c,al_ac1e65eb[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5aeea78d (
    .a(al_5e11d7be[18]),
    .b(al_6d689829[18]),
    .c(al_e55eeb92),
    .o({al_2bd76071,al_ac1e65eb[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88e7db74 (
    .a(al_5e11d7be[19]),
    .b(al_6d689829[19]),
    .c(al_2bd76071),
    .o({al_f5c68653,al_ac1e65eb[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9286c06e (
    .a(al_5e11d7be[20]),
    .b(al_6d689829[20]),
    .c(al_f5c68653),
    .o({al_7b6818a7,al_ac1e65eb[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ea9ec98 (
    .a(al_5e11d7be[21]),
    .b(al_6d689829[21]),
    .c(al_7b6818a7),
    .o({al_ce1229f8,al_ac1e65eb[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b6df570d (
    .a(al_5e11d7be[22]),
    .b(al_6d689829[22]),
    .c(al_ce1229f8),
    .o({al_77221701,al_ac1e65eb[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b2fe22e7 (
    .a(al_5e11d7be[23]),
    .b(al_6d689829[23]),
    .c(al_77221701),
    .o({al_c6a9c727,al_ac1e65eb[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bca11881 (
    .a(al_5e11d7be[24]),
    .b(al_6d689829[24]),
    .c(al_c6a9c727),
    .o({al_e5f7a519,al_ac1e65eb[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b7e3955 (
    .a(al_5e11d7be[25]),
    .b(al_6d689829[25]),
    .c(al_e5f7a519),
    .o({al_c65e25f4,al_ac1e65eb[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d82e5cce (
    .a(al_5e11d7be[26]),
    .b(al_6d689829[26]),
    .c(al_c65e25f4),
    .o({al_a839234c,al_ac1e65eb[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5fd41b50 (
    .a(al_5e11d7be[27]),
    .b(al_6d689829[27]),
    .c(al_a839234c),
    .o({al_e0116105,al_ac1e65eb[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8334f2d1 (
    .a(al_5e11d7be[1]),
    .b(al_6d689829[1]),
    .c(al_4b7e6f4c),
    .o({al_dc48d934,al_ac1e65eb[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_165a4d71 (
    .a(al_5e11d7be[28]),
    .b(al_6d689829[28]),
    .c(al_e0116105),
    .o({open_n35,al_ac1e65eb[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa68e50a (
    .a(al_5e11d7be[2]),
    .b(al_6d689829[2]),
    .c(al_dc48d934),
    .o({al_65f78d31,al_ac1e65eb[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f535854f (
    .a(al_5e11d7be[3]),
    .b(al_6d689829[3]),
    .c(al_65f78d31),
    .o({al_9f58115d,al_ac1e65eb[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47acf8fd (
    .a(al_5e11d7be[4]),
    .b(al_6d689829[4]),
    .c(al_9f58115d),
    .o({al_6678a2d9,al_ac1e65eb[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfff5f88 (
    .a(al_5e11d7be[5]),
    .b(al_6d689829[5]),
    .c(al_6678a2d9),
    .o({al_d662cc5f,al_ac1e65eb[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5dc05aa (
    .a(al_5e11d7be[6]),
    .b(al_6d689829[6]),
    .c(al_d662cc5f),
    .o({al_121b0ac0,al_ac1e65eb[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc4ce8ed (
    .a(al_5e11d7be[7]),
    .b(al_6d689829[7]),
    .c(al_121b0ac0),
    .o({al_74c02a6e,al_ac1e65eb[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_31460b8a (
    .a(1'b0),
    .o({al_b7706566,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a40d1df8 (
    .a(al_2c916a43[8]),
    .b(al_62f4aab[8]),
    .c(al_a8099213),
    .o({al_89797e8b,al_4e1fa175[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_64b8b6e8 (
    .a(al_2c916a43[9]),
    .b(al_62f4aab[9]),
    .c(al_89797e8b),
    .o({al_d4fb750d,al_4e1fa175[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98a55e98 (
    .a(al_2c916a43[10]),
    .b(al_62f4aab[10]),
    .c(al_d4fb750d),
    .o({al_c0a4beaf,al_4e1fa175[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a91b1aa (
    .a(al_2c916a43[11]),
    .b(al_62f4aab[11]),
    .c(al_c0a4beaf),
    .o({al_f1885c7b,al_4e1fa175[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3cde8b3d (
    .a(al_2c916a43[12]),
    .b(al_62f4aab[12]),
    .c(al_f1885c7b),
    .o({al_406fb43d,al_4e1fa175[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_77103919 (
    .a(al_2c916a43[13]),
    .b(al_62f4aab[13]),
    .c(al_406fb43d),
    .o({al_2ae006a6,al_4e1fa175[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b13a6286 (
    .a(al_2c916a43[14]),
    .b(al_62f4aab[14]),
    .c(al_2ae006a6),
    .o({al_25a1ab81,al_4e1fa175[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ed28c8d (
    .a(al_2c916a43[15]),
    .b(al_62f4aab[15]),
    .c(al_25a1ab81),
    .o({al_7bc6bbc7,al_4e1fa175[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2278d9d1 (
    .a(al_2c916a43[16]),
    .b(al_62f4aab[16]),
    .c(al_7bc6bbc7),
    .o({al_5d510d59,al_4e1fa175[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a953d37d (
    .a(al_2c916a43[17]),
    .b(al_62f4aab[17]),
    .c(al_5d510d59),
    .o({al_d82381d,al_4e1fa175[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d4bdeed7 (
    .a(al_2c916a43[0]),
    .b(al_62f4aab[0]),
    .c(al_b7706566),
    .o({al_32713696,al_4e1fa175[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_815ddabb (
    .a(al_2c916a43[18]),
    .b(al_62f4aab[18]),
    .c(al_d82381d),
    .o({al_9f37eb9f,al_4e1fa175[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c765fcf2 (
    .a(al_2c916a43[19]),
    .b(al_62f4aab[19]),
    .c(al_9f37eb9f),
    .o({al_3fca7,al_4e1fa175[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_998edeed (
    .a(al_2c916a43[20]),
    .b(al_62f4aab[20]),
    .c(al_3fca7),
    .o({al_22c2b9e6,al_4e1fa175[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ac02da8 (
    .a(al_2c916a43[21]),
    .b(al_62f4aab[21]),
    .c(al_22c2b9e6),
    .o({al_72694321,al_4e1fa175[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8c41e823 (
    .a(al_2c916a43[22]),
    .b(al_62f4aab[22]),
    .c(al_72694321),
    .o({al_5e0efc9d,al_4e1fa175[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d1a9f60a (
    .a(al_2c916a43[23]),
    .b(al_62f4aab[23]),
    .c(al_5e0efc9d),
    .o({al_4218870a,al_4e1fa175[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c57e73d (
    .a(al_2c916a43[24]),
    .b(al_62f4aab[24]),
    .c(al_4218870a),
    .o({al_debafe7e,al_4e1fa175[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b43bab3f (
    .a(al_2c916a43[25]),
    .b(al_62f4aab[25]),
    .c(al_debafe7e),
    .o({al_fd1c7e35,al_4e1fa175[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88448bc9 (
    .a(al_2c916a43[26]),
    .b(al_62f4aab[26]),
    .c(al_fd1c7e35),
    .o({al_f4a4c863,al_4e1fa175[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce4ca9e0 (
    .a(al_2c916a43[27]),
    .b(al_62f4aab[27]),
    .c(al_f4a4c863),
    .o({al_47aec73d,al_4e1fa175[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5e23e14 (
    .a(al_2c916a43[1]),
    .b(al_62f4aab[1]),
    .c(al_32713696),
    .o({al_58c1d211,al_4e1fa175[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c0758015 (
    .a(al_2c916a43[28]),
    .b(al_62f4aab[28]),
    .c(al_47aec73d),
    .o({open_n39,al_4e1fa175[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd207d59 (
    .a(al_2c916a43[2]),
    .b(al_62f4aab[2]),
    .c(al_58c1d211),
    .o({al_f6e6833c,al_4e1fa175[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_465c7c96 (
    .a(al_2c916a43[3]),
    .b(al_62f4aab[3]),
    .c(al_f6e6833c),
    .o({al_d6b08360,al_4e1fa175[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b997726c (
    .a(al_2c916a43[4]),
    .b(al_62f4aab[4]),
    .c(al_d6b08360),
    .o({al_ab39c04d,al_4e1fa175[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8cc46a2 (
    .a(al_2c916a43[5]),
    .b(al_62f4aab[5]),
    .c(al_ab39c04d),
    .o({al_a1a76be0,al_4e1fa175[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_85fbc719 (
    .a(al_2c916a43[6]),
    .b(al_62f4aab[6]),
    .c(al_a1a76be0),
    .o({al_80b80f4,al_4e1fa175[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c7a2c613 (
    .a(al_2c916a43[7]),
    .b(al_62f4aab[7]),
    .c(al_80b80f4),
    .o({al_a8099213,al_4e1fa175[7]}));

endmodule 

